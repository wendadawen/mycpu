`timescale 1ns / 1ps


module mips(
	input wire clk,rst,
	output wire[31:0] pcF,
	input wire[31:0] instrF,
	output wire memwriteM,
	output wire[31:0] aluoutM,writedataM,
	input wire[31:0] readdataM
);
	
	wire [5:0] opD,functD;
	wire regdstE,alusrcE,pcsrcD,jumpD;
	wire [1:0] memtoregE,memtoregM,memtoregW;
	wire regwriteE,regwriteM,regwriteW;
	wire [7:0] alucontrolE;
	wire LoWrite_E, HiWrite_E;
	wire LoSrc_E, HiSrc_E;
	wire flushE,equalD;
	wire Stall_E, Flush_M;

	controller c(
		clk,rst,
		//decode stage
		opD,functD,equalD,
		pcsrcD,branchD,jumpD,
		
		//execute stage
		flushE,
		memtoregE,alusrcE,
		regdstE,regwriteE,	
		alucontrolE,
		LoWrite_E, HiWrite_E,
		LoSrc_E, HiSrc_E,
		Stall_E,

		//mem stage
		memtoregM,memwriteM,
		regwriteM,
		Flush_M,

		//write back stage
		memtoregW,regwriteW
	);
	datapath dp(
		clk,rst,
		//fetch stage
		pcF,
		instrF,
		//decode stage
		pcsrcD,branchD,
		jumpD,
		equalD,
		opD,functD,
		//execute stage
		memtoregE,
		alusrcE,regdstE,
		regwriteE,
		alucontrolE,
		flushE,
		LoWrite_E, HiWrite_E,
		LoSrc_E, HiSrc_E,
		Stall_E,
		//mem stage
		memtoregM,
		regwriteM,
		aluoutM,writedataM,
		readdataM,
		Flush_M,
		//writeback stage
		memtoregW,
		regwriteW
	);
	
endmodule
